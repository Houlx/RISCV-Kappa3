module vector_reg(input clock,
                    input reset,
                    
                    input [4:0] vs1_addr,
                    input [4:0] vs2_addr,
                    input [4:0] vd_addr,

                    input [] in,
                    input ld,

                    output [] vs1_out,
                    output [] vs2_out
                    );
endmodule